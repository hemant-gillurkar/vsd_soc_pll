magic
tech sky130A
magscale 1 2
timestamp 1613927320
<< obsli1 >>
rect 44 113814 717556 924551
<< obsm1 >>
rect 0 47812 717600 990276
<< obsm2 >>
rect 0 47806 717600 990282
<< obsm3 >>
rect 0 113648 717600 924540
<< obsm4 >>
rect 0 0 717600 1037600
<< metal5 >>
rect 1152 1032681 716448 1033001
rect 1152 1017363 716448 1017683
rect 1152 1002045 716448 1002365
rect 1152 986727 716448 987047
rect 1152 971409 716448 971729
rect 1152 956091 716448 956411
rect 1152 940773 716448 941093
rect 1152 925455 716448 925775
rect 1152 910137 716448 910457
rect 1152 894819 716448 895139
rect 1152 879501 716448 879821
rect 1152 864183 716448 864503
rect 1152 848865 716448 849185
rect 1152 833547 716448 833867
rect 1152 818229 716448 818549
rect 1152 802911 716448 803231
rect 1152 787593 716448 787913
rect 1152 772275 716448 772595
rect 1152 756957 716448 757277
rect 1152 741639 716448 741959
rect 1152 726321 716448 726641
rect 1152 711003 716448 711323
rect 1152 695685 716448 696005
rect 1152 680367 716448 680687
rect 1152 665049 716448 665369
rect 1152 649731 716448 650051
rect 1152 634413 716448 634733
rect 1152 619095 716448 619415
rect 1152 603777 716448 604097
rect 1152 588459 716448 588779
rect 1152 573141 716448 573461
rect 1152 557823 716448 558143
rect 1152 542505 716448 542825
rect 1152 527187 716448 527507
rect 1152 511869 716448 512189
rect 1152 496551 716448 496871
rect 1152 481233 716448 481553
rect 1152 465915 716448 466235
rect 1152 450597 716448 450917
rect 1152 435279 716448 435599
rect 1152 419961 716448 420281
rect 1152 404643 716448 404963
rect 1152 389325 716448 389645
rect 1152 374007 716448 374327
rect 1152 358689 716448 359009
rect 1152 343371 716448 343691
rect 1152 328053 716448 328373
rect 1152 312735 716448 313055
rect 1152 297417 716448 297737
rect 1152 282099 716448 282419
rect 1152 266781 716448 267101
rect 1152 251463 716448 251783
rect 1152 236145 716448 236465
rect 1152 220827 716448 221147
rect 1152 205509 716448 205829
rect 1152 190191 716448 190511
rect 1152 174873 716448 175193
rect 1152 159555 716448 159875
rect 1152 144237 716448 144557
rect 1152 128919 716448 129239
rect 1152 113601 716448 113921
rect 1152 98283 716448 98603
rect 1152 82965 716448 83285
rect 1152 67647 716448 67967
rect 1152 52329 716448 52649
rect 1152 37011 716448 37331
rect 1152 21693 716448 22013
rect 1152 6375 716448 6695
<< obsm5 >>
rect 0 1033321 717600 1037600
rect 0 1032361 832 1033321
rect 716768 1032361 717600 1033321
rect 0 1018003 717600 1032361
rect 0 1017043 832 1018003
rect 716768 1017043 717600 1018003
rect 0 1002685 717600 1017043
rect 0 1001725 832 1002685
rect 716768 1001725 717600 1002685
rect 0 987367 717600 1001725
rect 0 986407 832 987367
rect 716768 986407 717600 987367
rect 0 972049 717600 986407
rect 0 971089 832 972049
rect 716768 971089 717600 972049
rect 0 956731 717600 971089
rect 0 955771 832 956731
rect 716768 955771 717600 956731
rect 0 941413 717600 955771
rect 0 940453 832 941413
rect 716768 940453 717600 941413
rect 0 926095 717600 940453
rect 0 925135 832 926095
rect 716768 925135 717600 926095
rect 0 910777 717600 925135
rect 0 909817 832 910777
rect 716768 909817 717600 910777
rect 0 895459 717600 909817
rect 0 894499 832 895459
rect 716768 894499 717600 895459
rect 0 880141 717600 894499
rect 0 879181 832 880141
rect 716768 879181 717600 880141
rect 0 864823 717600 879181
rect 0 863863 832 864823
rect 716768 863863 717600 864823
rect 0 849505 717600 863863
rect 0 848545 832 849505
rect 716768 848545 717600 849505
rect 0 834187 717600 848545
rect 0 833227 832 834187
rect 716768 833227 717600 834187
rect 0 818869 717600 833227
rect 0 817909 832 818869
rect 716768 817909 717600 818869
rect 0 803551 717600 817909
rect 0 802591 832 803551
rect 716768 802591 717600 803551
rect 0 788233 717600 802591
rect 0 787273 832 788233
rect 716768 787273 717600 788233
rect 0 772915 717600 787273
rect 0 771955 832 772915
rect 716768 771955 717600 772915
rect 0 757597 717600 771955
rect 0 756637 832 757597
rect 716768 756637 717600 757597
rect 0 742279 717600 756637
rect 0 741319 832 742279
rect 716768 741319 717600 742279
rect 0 726961 717600 741319
rect 0 726001 832 726961
rect 716768 726001 717600 726961
rect 0 711643 717600 726001
rect 0 710683 832 711643
rect 716768 710683 717600 711643
rect 0 696325 717600 710683
rect 0 695365 832 696325
rect 716768 695365 717600 696325
rect 0 681007 717600 695365
rect 0 680047 832 681007
rect 716768 680047 717600 681007
rect 0 665689 717600 680047
rect 0 664729 832 665689
rect 716768 664729 717600 665689
rect 0 650371 717600 664729
rect 0 649411 832 650371
rect 716768 649411 717600 650371
rect 0 635053 717600 649411
rect 0 634093 832 635053
rect 716768 634093 717600 635053
rect 0 619735 717600 634093
rect 0 618775 832 619735
rect 716768 618775 717600 619735
rect 0 604417 717600 618775
rect 0 603457 832 604417
rect 716768 603457 717600 604417
rect 0 589099 717600 603457
rect 0 588139 832 589099
rect 716768 588139 717600 589099
rect 0 573781 717600 588139
rect 0 572821 832 573781
rect 716768 572821 717600 573781
rect 0 558463 717600 572821
rect 0 557503 832 558463
rect 716768 557503 717600 558463
rect 0 543145 717600 557503
rect 0 542185 832 543145
rect 716768 542185 717600 543145
rect 0 527827 717600 542185
rect 0 526867 832 527827
rect 716768 526867 717600 527827
rect 0 512509 717600 526867
rect 0 511549 832 512509
rect 716768 511549 717600 512509
rect 0 497191 717600 511549
rect 0 496231 832 497191
rect 716768 496231 717600 497191
rect 0 481873 717600 496231
rect 0 480913 832 481873
rect 716768 480913 717600 481873
rect 0 466555 717600 480913
rect 0 465595 832 466555
rect 716768 465595 717600 466555
rect 0 451237 717600 465595
rect 0 450277 832 451237
rect 716768 450277 717600 451237
rect 0 435919 717600 450277
rect 0 434959 832 435919
rect 716768 434959 717600 435919
rect 0 420601 717600 434959
rect 0 419641 832 420601
rect 716768 419641 717600 420601
rect 0 405283 717600 419641
rect 0 404323 832 405283
rect 716768 404323 717600 405283
rect 0 389965 717600 404323
rect 0 389005 832 389965
rect 716768 389005 717600 389965
rect 0 374647 717600 389005
rect 0 373687 832 374647
rect 716768 373687 717600 374647
rect 0 359329 717600 373687
rect 0 358369 832 359329
rect 716768 358369 717600 359329
rect 0 344011 717600 358369
rect 0 343051 832 344011
rect 716768 343051 717600 344011
rect 0 328693 717600 343051
rect 0 327733 832 328693
rect 716768 327733 717600 328693
rect 0 313375 717600 327733
rect 0 312415 832 313375
rect 716768 312415 717600 313375
rect 0 298057 717600 312415
rect 0 297097 832 298057
rect 716768 297097 717600 298057
rect 0 282739 717600 297097
rect 0 281779 832 282739
rect 716768 281779 717600 282739
rect 0 267421 717600 281779
rect 0 266461 832 267421
rect 716768 266461 717600 267421
rect 0 252103 717600 266461
rect 0 251143 832 252103
rect 716768 251143 717600 252103
rect 0 236785 717600 251143
rect 0 235825 832 236785
rect 716768 235825 717600 236785
rect 0 221467 717600 235825
rect 0 220507 832 221467
rect 716768 220507 717600 221467
rect 0 206149 717600 220507
rect 0 205189 832 206149
rect 716768 205189 717600 206149
rect 0 190831 717600 205189
rect 0 189871 832 190831
rect 716768 189871 717600 190831
rect 0 175513 717600 189871
rect 0 174553 832 175513
rect 716768 174553 717600 175513
rect 0 160195 717600 174553
rect 0 159235 832 160195
rect 716768 159235 717600 160195
rect 0 144877 717600 159235
rect 0 143917 832 144877
rect 716768 143917 717600 144877
rect 0 129559 717600 143917
rect 0 128599 832 129559
rect 716768 128599 717600 129559
rect 0 114241 717600 128599
rect 0 113281 832 114241
rect 716768 113281 717600 114241
rect 0 98923 717600 113281
rect 0 97963 832 98923
rect 716768 97963 717600 98923
rect 0 83605 717600 97963
rect 0 82645 832 83605
rect 716768 82645 717600 83605
rect 0 68287 717600 82645
rect 0 67327 832 68287
rect 716768 67327 717600 68287
rect 0 52969 717600 67327
rect 0 52009 832 52969
rect 716768 52009 717600 52969
rect 0 37651 717600 52009
rect 0 36691 832 37651
rect 716768 36691 717600 37651
rect 0 22333 717600 36691
rect 0 21373 832 22333
rect 716768 21373 717600 22333
rect 0 7015 717600 21373
rect 0 6055 832 7015
rect 716768 6055 717600 7015
rect 0 0 717600 6055
<< labels >>
rlabel metal5 s 1152 1017363 716448 1017683 6 VPWR
port 1 nsew power bidirectional
rlabel metal5 s 1152 986727 716448 987047 6 VPWR.extra1
port 2 nsew power bidirectional
rlabel metal5 s 1152 956091 716448 956411 6 VPWR.extra2
port 3 nsew power bidirectional
rlabel metal5 s 1152 925455 716448 925775 6 VPWR.extra3
port 4 nsew power bidirectional
rlabel metal5 s 1152 894819 716448 895139 6 VPWR.extra4
port 5 nsew power bidirectional
rlabel metal5 s 1152 864183 716448 864503 6 VPWR.extra5
port 6 nsew power bidirectional
rlabel metal5 s 1152 833547 716448 833867 6 VPWR.extra6
port 7 nsew power bidirectional
rlabel metal5 s 1152 802911 716448 803231 6 VPWR.extra7
port 8 nsew power bidirectional
rlabel metal5 s 1152 772275 716448 772595 6 VPWR.extra8
port 9 nsew power bidirectional
rlabel metal5 s 1152 741639 716448 741959 6 VPWR.extra9
port 10 nsew power bidirectional
rlabel metal5 s 1152 711003 716448 711323 6 VPWR.extra10
port 11 nsew power bidirectional
rlabel metal5 s 1152 680367 716448 680687 6 VPWR.extra11
port 12 nsew power bidirectional
rlabel metal5 s 1152 649731 716448 650051 6 VPWR.extra12
port 13 nsew power bidirectional
rlabel metal5 s 1152 619095 716448 619415 6 VPWR.extra13
port 14 nsew power bidirectional
rlabel metal5 s 1152 588459 716448 588779 6 VPWR.extra14
port 15 nsew power bidirectional
rlabel metal5 s 1152 557823 716448 558143 6 VPWR.extra15
port 16 nsew power bidirectional
rlabel metal5 s 1152 527187 716448 527507 6 VPWR.extra16
port 17 nsew power bidirectional
rlabel metal5 s 1152 496551 716448 496871 6 VPWR.extra17
port 18 nsew power bidirectional
rlabel metal5 s 1152 465915 716448 466235 6 VPWR.extra18
port 19 nsew power bidirectional
rlabel metal5 s 1152 435279 716448 435599 6 VPWR.extra19
port 20 nsew power bidirectional
rlabel metal5 s 1152 404643 716448 404963 6 VPWR.extra20
port 21 nsew power bidirectional
rlabel metal5 s 1152 374007 716448 374327 6 VPWR.extra21
port 22 nsew power bidirectional
rlabel metal5 s 1152 343371 716448 343691 6 VPWR.extra22
port 23 nsew power bidirectional
rlabel metal5 s 1152 312735 716448 313055 6 VPWR.extra23
port 24 nsew power bidirectional
rlabel metal5 s 1152 282099 716448 282419 6 VPWR.extra24
port 25 nsew power bidirectional
rlabel metal5 s 1152 251463 716448 251783 6 VPWR.extra25
port 26 nsew power bidirectional
rlabel metal5 s 1152 220827 716448 221147 6 VPWR.extra26
port 27 nsew power bidirectional
rlabel metal5 s 1152 190191 716448 190511 6 VPWR.extra27
port 28 nsew power bidirectional
rlabel metal5 s 1152 159555 716448 159875 6 VPWR.extra28
port 29 nsew power bidirectional
rlabel metal5 s 1152 128919 716448 129239 6 VPWR.extra29
port 30 nsew power bidirectional
rlabel metal5 s 1152 98283 716448 98603 6 VPWR.extra30
port 31 nsew power bidirectional
rlabel metal5 s 1152 67647 716448 67967 6 VPWR.extra31
port 32 nsew power bidirectional
rlabel metal5 s 1152 37011 716448 37331 6 VPWR.extra32
port 33 nsew power bidirectional
rlabel metal5 s 1152 6375 716448 6695 6 VPWR.extra33
port 34 nsew power bidirectional
rlabel metal5 s 1152 1032681 716448 1033001 6 VGND
port 35 nsew ground bidirectional
rlabel metal5 s 1152 1002045 716448 1002365 6 VGND.extra1
port 36 nsew ground bidirectional
rlabel metal5 s 1152 971409 716448 971729 6 VGND.extra2
port 37 nsew ground bidirectional
rlabel metal5 s 1152 940773 716448 941093 6 VGND.extra3
port 38 nsew ground bidirectional
rlabel metal5 s 1152 910137 716448 910457 6 VGND.extra4
port 39 nsew ground bidirectional
rlabel metal5 s 1152 879501 716448 879821 6 VGND.extra5
port 40 nsew ground bidirectional
rlabel metal5 s 1152 848865 716448 849185 6 VGND.extra6
port 41 nsew ground bidirectional
rlabel metal5 s 1152 818229 716448 818549 6 VGND.extra7
port 42 nsew ground bidirectional
rlabel metal5 s 1152 787593 716448 787913 6 VGND.extra8
port 43 nsew ground bidirectional
rlabel metal5 s 1152 756957 716448 757277 6 VGND.extra9
port 44 nsew ground bidirectional
rlabel metal5 s 1152 726321 716448 726641 6 VGND.extra10
port 45 nsew ground bidirectional
rlabel metal5 s 1152 695685 716448 696005 6 VGND.extra11
port 46 nsew ground bidirectional
rlabel metal5 s 1152 665049 716448 665369 6 VGND.extra12
port 47 nsew ground bidirectional
rlabel metal5 s 1152 634413 716448 634733 6 VGND.extra13
port 48 nsew ground bidirectional
rlabel metal5 s 1152 603777 716448 604097 6 VGND.extra14
port 49 nsew ground bidirectional
rlabel metal5 s 1152 573141 716448 573461 6 VGND.extra15
port 50 nsew ground bidirectional
rlabel metal5 s 1152 542505 716448 542825 6 VGND.extra16
port 51 nsew ground bidirectional
rlabel metal5 s 1152 511869 716448 512189 6 VGND.extra17
port 52 nsew ground bidirectional
rlabel metal5 s 1152 481233 716448 481553 6 VGND.extra18
port 53 nsew ground bidirectional
rlabel metal5 s 1152 450597 716448 450917 6 VGND.extra19
port 54 nsew ground bidirectional
rlabel metal5 s 1152 419961 716448 420281 6 VGND.extra20
port 55 nsew ground bidirectional
rlabel metal5 s 1152 389325 716448 389645 6 VGND.extra21
port 56 nsew ground bidirectional
rlabel metal5 s 1152 358689 716448 359009 6 VGND.extra22
port 57 nsew ground bidirectional
rlabel metal5 s 1152 328053 716448 328373 6 VGND.extra23
port 58 nsew ground bidirectional
rlabel metal5 s 1152 297417 716448 297737 6 VGND.extra24
port 59 nsew ground bidirectional
rlabel metal5 s 1152 266781 716448 267101 6 VGND.extra25
port 60 nsew ground bidirectional
rlabel metal5 s 1152 236145 716448 236465 6 VGND.extra26
port 61 nsew ground bidirectional
rlabel metal5 s 1152 205509 716448 205829 6 VGND.extra27
port 62 nsew ground bidirectional
rlabel metal5 s 1152 174873 716448 175193 6 VGND.extra28
port 63 nsew ground bidirectional
rlabel metal5 s 1152 144237 716448 144557 6 VGND.extra29
port 64 nsew ground bidirectional
rlabel metal5 s 1152 113601 716448 113921 6 VGND.extra30
port 65 nsew ground bidirectional
rlabel metal5 s 1152 82965 716448 83285 6 VGND.extra31
port 66 nsew ground bidirectional
rlabel metal5 s 1152 52329 716448 52649 6 VGND.extra32
port 67 nsew ground bidirectional
rlabel metal5 s 1152 21693 716448 22013 6 VGND.extra33
port 68 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 717600 1037600
string LEFview TRUE
<< end >>
