VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO vsdPLLSoC
  CLASS BLOCK ;
  FOREIGN vsdPLLSoC ;
  ORIGIN 0.000 0.000 ;
  SIZE 3588.000 BY 5188.000 ;
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.760 5086.815 3582.240 5088.415 ;
    END
  END VPWR
  PIN VPWR.extra1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.760 4933.635 3582.240 4935.235 ;
    END
  END VPWR.extra1
  PIN VPWR.extra2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.760 4780.455 3582.240 4782.055 ;
    END
  END VPWR.extra2
  PIN VPWR.extra3
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.760 4627.275 3582.240 4628.875 ;
    END
  END VPWR.extra3
  PIN VPWR.extra4
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.760 4474.095 3582.240 4475.695 ;
    END
  END VPWR.extra4
  PIN VPWR.extra5
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.760 4320.915 3582.240 4322.515 ;
    END
  END VPWR.extra5
  PIN VPWR.extra6
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.760 4167.735 3582.240 4169.335 ;
    END
  END VPWR.extra6
  PIN VPWR.extra7
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.760 4014.555 3582.240 4016.155 ;
    END
  END VPWR.extra7
  PIN VPWR.extra8
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.760 3861.375 3582.240 3862.975 ;
    END
  END VPWR.extra8
  PIN VPWR.extra9
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.760 3708.195 3582.240 3709.795 ;
    END
  END VPWR.extra9
  PIN VPWR.extra10
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.760 3555.015 3582.240 3556.615 ;
    END
  END VPWR.extra10
  PIN VPWR.extra11
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.760 3401.835 3582.240 3403.435 ;
    END
  END VPWR.extra11
  PIN VPWR.extra12
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.760 3248.655 3582.240 3250.255 ;
    END
  END VPWR.extra12
  PIN VPWR.extra13
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.760 3095.475 3582.240 3097.075 ;
    END
  END VPWR.extra13
  PIN VPWR.extra14
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.760 2942.295 3582.240 2943.895 ;
    END
  END VPWR.extra14
  PIN VPWR.extra15
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.760 2789.115 3582.240 2790.715 ;
    END
  END VPWR.extra15
  PIN VPWR.extra16
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.760 2635.935 3582.240 2637.535 ;
    END
  END VPWR.extra16
  PIN VPWR.extra17
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.760 2482.755 3582.240 2484.355 ;
    END
  END VPWR.extra17
  PIN VPWR.extra18
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.760 2329.575 3582.240 2331.175 ;
    END
  END VPWR.extra18
  PIN VPWR.extra19
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.760 2176.395 3582.240 2177.995 ;
    END
  END VPWR.extra19
  PIN VPWR.extra20
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.760 2023.215 3582.240 2024.815 ;
    END
  END VPWR.extra20
  PIN VPWR.extra21
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.760 1870.035 3582.240 1871.635 ;
    END
  END VPWR.extra21
  PIN VPWR.extra22
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.760 1716.855 3582.240 1718.455 ;
    END
  END VPWR.extra22
  PIN VPWR.extra23
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.760 1563.675 3582.240 1565.275 ;
    END
  END VPWR.extra23
  PIN VPWR.extra24
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.760 1410.495 3582.240 1412.095 ;
    END
  END VPWR.extra24
  PIN VPWR.extra25
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.760 1257.315 3582.240 1258.915 ;
    END
  END VPWR.extra25
  PIN VPWR.extra26
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.760 1104.135 3582.240 1105.735 ;
    END
  END VPWR.extra26
  PIN VPWR.extra27
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.760 950.955 3582.240 952.555 ;
    END
  END VPWR.extra27
  PIN VPWR.extra28
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.760 797.775 3582.240 799.375 ;
    END
  END VPWR.extra28
  PIN VPWR.extra29
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.760 644.595 3582.240 646.195 ;
    END
  END VPWR.extra29
  PIN VPWR.extra30
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.760 491.415 3582.240 493.015 ;
    END
  END VPWR.extra30
  PIN VPWR.extra31
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.760 338.235 3582.240 339.835 ;
    END
  END VPWR.extra31
  PIN VPWR.extra32
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.760 185.055 3582.240 186.655 ;
    END
  END VPWR.extra32
  PIN VPWR.extra33
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.760 31.875 3582.240 33.475 ;
    END
  END VPWR.extra33
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.760 5163.405 3582.240 5165.005 ;
    END
  END VGND
  PIN VGND.extra1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.760 5010.225 3582.240 5011.825 ;
    END
  END VGND.extra1
  PIN VGND.extra2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.760 4857.045 3582.240 4858.645 ;
    END
  END VGND.extra2
  PIN VGND.extra3
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.760 4703.865 3582.240 4705.465 ;
    END
  END VGND.extra3
  PIN VGND.extra4
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.760 4550.685 3582.240 4552.285 ;
    END
  END VGND.extra4
  PIN VGND.extra5
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.760 4397.505 3582.240 4399.105 ;
    END
  END VGND.extra5
  PIN VGND.extra6
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.760 4244.325 3582.240 4245.925 ;
    END
  END VGND.extra6
  PIN VGND.extra7
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.760 4091.145 3582.240 4092.745 ;
    END
  END VGND.extra7
  PIN VGND.extra8
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.760 3937.965 3582.240 3939.565 ;
    END
  END VGND.extra8
  PIN VGND.extra9
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.760 3784.785 3582.240 3786.385 ;
    END
  END VGND.extra9
  PIN VGND.extra10
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.760 3631.605 3582.240 3633.205 ;
    END
  END VGND.extra10
  PIN VGND.extra11
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.760 3478.425 3582.240 3480.025 ;
    END
  END VGND.extra11
  PIN VGND.extra12
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.760 3325.245 3582.240 3326.845 ;
    END
  END VGND.extra12
  PIN VGND.extra13
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.760 3172.065 3582.240 3173.665 ;
    END
  END VGND.extra13
  PIN VGND.extra14
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.760 3018.885 3582.240 3020.485 ;
    END
  END VGND.extra14
  PIN VGND.extra15
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.760 2865.705 3582.240 2867.305 ;
    END
  END VGND.extra15
  PIN VGND.extra16
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.760 2712.525 3582.240 2714.125 ;
    END
  END VGND.extra16
  PIN VGND.extra17
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.760 2559.345 3582.240 2560.945 ;
    END
  END VGND.extra17
  PIN VGND.extra18
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.760 2406.165 3582.240 2407.765 ;
    END
  END VGND.extra18
  PIN VGND.extra19
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.760 2252.985 3582.240 2254.585 ;
    END
  END VGND.extra19
  PIN VGND.extra20
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.760 2099.805 3582.240 2101.405 ;
    END
  END VGND.extra20
  PIN VGND.extra21
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.760 1946.625 3582.240 1948.225 ;
    END
  END VGND.extra21
  PIN VGND.extra22
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.760 1793.445 3582.240 1795.045 ;
    END
  END VGND.extra22
  PIN VGND.extra23
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.760 1640.265 3582.240 1641.865 ;
    END
  END VGND.extra23
  PIN VGND.extra24
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.760 1487.085 3582.240 1488.685 ;
    END
  END VGND.extra24
  PIN VGND.extra25
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.760 1333.905 3582.240 1335.505 ;
    END
  END VGND.extra25
  PIN VGND.extra26
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.760 1180.725 3582.240 1182.325 ;
    END
  END VGND.extra26
  PIN VGND.extra27
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.760 1027.545 3582.240 1029.145 ;
    END
  END VGND.extra27
  PIN VGND.extra28
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.760 874.365 3582.240 875.965 ;
    END
  END VGND.extra28
  PIN VGND.extra29
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.760 721.185 3582.240 722.785 ;
    END
  END VGND.extra29
  PIN VGND.extra30
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.760 568.005 3582.240 569.605 ;
    END
  END VGND.extra30
  PIN VGND.extra31
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.760 414.825 3582.240 416.425 ;
    END
  END VGND.extra31
  PIN VGND.extra32
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.760 261.645 3582.240 263.245 ;
    END
  END VGND.extra32
  PIN VGND.extra33
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.760 108.465 3582.240 110.065 ;
    END
  END VGND.extra33
  OBS
      LAYER li1 ;
        RECT 0.220 569.070 3587.780 4622.755 ;
      LAYER met1 ;
        RECT 0.000 239.060 3588.000 4951.380 ;
      LAYER met2 ;
        RECT 0.000 239.030 3588.000 4951.410 ;
      LAYER met3 ;
        RECT 0.000 568.240 3588.000 4622.700 ;
      LAYER met4 ;
        RECT 0.000 0.000 3588.000 5188.000 ;
      LAYER met5 ;
        RECT 0.000 5166.605 3588.000 5188.000 ;
        RECT 0.000 5161.805 4.160 5166.605 ;
        RECT 3583.840 5161.805 3588.000 5166.605 ;
        RECT 0.000 5090.015 3588.000 5161.805 ;
        RECT 0.000 5085.215 4.160 5090.015 ;
        RECT 3583.840 5085.215 3588.000 5090.015 ;
        RECT 0.000 5013.425 3588.000 5085.215 ;
        RECT 0.000 5008.625 4.160 5013.425 ;
        RECT 3583.840 5008.625 3588.000 5013.425 ;
        RECT 0.000 4936.835 3588.000 5008.625 ;
        RECT 0.000 4932.035 4.160 4936.835 ;
        RECT 3583.840 4932.035 3588.000 4936.835 ;
        RECT 0.000 4860.245 3588.000 4932.035 ;
        RECT 0.000 4855.445 4.160 4860.245 ;
        RECT 3583.840 4855.445 3588.000 4860.245 ;
        RECT 0.000 4783.655 3588.000 4855.445 ;
        RECT 0.000 4778.855 4.160 4783.655 ;
        RECT 3583.840 4778.855 3588.000 4783.655 ;
        RECT 0.000 4707.065 3588.000 4778.855 ;
        RECT 0.000 4702.265 4.160 4707.065 ;
        RECT 3583.840 4702.265 3588.000 4707.065 ;
        RECT 0.000 4630.475 3588.000 4702.265 ;
        RECT 0.000 4625.675 4.160 4630.475 ;
        RECT 3583.840 4625.675 3588.000 4630.475 ;
        RECT 0.000 4553.885 3588.000 4625.675 ;
        RECT 0.000 4549.085 4.160 4553.885 ;
        RECT 3583.840 4549.085 3588.000 4553.885 ;
        RECT 0.000 4477.295 3588.000 4549.085 ;
        RECT 0.000 4472.495 4.160 4477.295 ;
        RECT 3583.840 4472.495 3588.000 4477.295 ;
        RECT 0.000 4400.705 3588.000 4472.495 ;
        RECT 0.000 4395.905 4.160 4400.705 ;
        RECT 3583.840 4395.905 3588.000 4400.705 ;
        RECT 0.000 4324.115 3588.000 4395.905 ;
        RECT 0.000 4319.315 4.160 4324.115 ;
        RECT 3583.840 4319.315 3588.000 4324.115 ;
        RECT 0.000 4247.525 3588.000 4319.315 ;
        RECT 0.000 4242.725 4.160 4247.525 ;
        RECT 3583.840 4242.725 3588.000 4247.525 ;
        RECT 0.000 4170.935 3588.000 4242.725 ;
        RECT 0.000 4166.135 4.160 4170.935 ;
        RECT 3583.840 4166.135 3588.000 4170.935 ;
        RECT 0.000 4094.345 3588.000 4166.135 ;
        RECT 0.000 4089.545 4.160 4094.345 ;
        RECT 3583.840 4089.545 3588.000 4094.345 ;
        RECT 0.000 4017.755 3588.000 4089.545 ;
        RECT 0.000 4012.955 4.160 4017.755 ;
        RECT 3583.840 4012.955 3588.000 4017.755 ;
        RECT 0.000 3941.165 3588.000 4012.955 ;
        RECT 0.000 3936.365 4.160 3941.165 ;
        RECT 3583.840 3936.365 3588.000 3941.165 ;
        RECT 0.000 3864.575 3588.000 3936.365 ;
        RECT 0.000 3859.775 4.160 3864.575 ;
        RECT 3583.840 3859.775 3588.000 3864.575 ;
        RECT 0.000 3787.985 3588.000 3859.775 ;
        RECT 0.000 3783.185 4.160 3787.985 ;
        RECT 3583.840 3783.185 3588.000 3787.985 ;
        RECT 0.000 3711.395 3588.000 3783.185 ;
        RECT 0.000 3706.595 4.160 3711.395 ;
        RECT 3583.840 3706.595 3588.000 3711.395 ;
        RECT 0.000 3634.805 3588.000 3706.595 ;
        RECT 0.000 3630.005 4.160 3634.805 ;
        RECT 3583.840 3630.005 3588.000 3634.805 ;
        RECT 0.000 3558.215 3588.000 3630.005 ;
        RECT 0.000 3553.415 4.160 3558.215 ;
        RECT 3583.840 3553.415 3588.000 3558.215 ;
        RECT 0.000 3481.625 3588.000 3553.415 ;
        RECT 0.000 3476.825 4.160 3481.625 ;
        RECT 3583.840 3476.825 3588.000 3481.625 ;
        RECT 0.000 3405.035 3588.000 3476.825 ;
        RECT 0.000 3400.235 4.160 3405.035 ;
        RECT 3583.840 3400.235 3588.000 3405.035 ;
        RECT 0.000 3328.445 3588.000 3400.235 ;
        RECT 0.000 3323.645 4.160 3328.445 ;
        RECT 3583.840 3323.645 3588.000 3328.445 ;
        RECT 0.000 3251.855 3588.000 3323.645 ;
        RECT 0.000 3247.055 4.160 3251.855 ;
        RECT 3583.840 3247.055 3588.000 3251.855 ;
        RECT 0.000 3175.265 3588.000 3247.055 ;
        RECT 0.000 3170.465 4.160 3175.265 ;
        RECT 3583.840 3170.465 3588.000 3175.265 ;
        RECT 0.000 3098.675 3588.000 3170.465 ;
        RECT 0.000 3093.875 4.160 3098.675 ;
        RECT 3583.840 3093.875 3588.000 3098.675 ;
        RECT 0.000 3022.085 3588.000 3093.875 ;
        RECT 0.000 3017.285 4.160 3022.085 ;
        RECT 3583.840 3017.285 3588.000 3022.085 ;
        RECT 0.000 2945.495 3588.000 3017.285 ;
        RECT 0.000 2940.695 4.160 2945.495 ;
        RECT 3583.840 2940.695 3588.000 2945.495 ;
        RECT 0.000 2868.905 3588.000 2940.695 ;
        RECT 0.000 2864.105 4.160 2868.905 ;
        RECT 3583.840 2864.105 3588.000 2868.905 ;
        RECT 0.000 2792.315 3588.000 2864.105 ;
        RECT 0.000 2787.515 4.160 2792.315 ;
        RECT 3583.840 2787.515 3588.000 2792.315 ;
        RECT 0.000 2715.725 3588.000 2787.515 ;
        RECT 0.000 2710.925 4.160 2715.725 ;
        RECT 3583.840 2710.925 3588.000 2715.725 ;
        RECT 0.000 2639.135 3588.000 2710.925 ;
        RECT 0.000 2634.335 4.160 2639.135 ;
        RECT 3583.840 2634.335 3588.000 2639.135 ;
        RECT 0.000 2562.545 3588.000 2634.335 ;
        RECT 0.000 2557.745 4.160 2562.545 ;
        RECT 3583.840 2557.745 3588.000 2562.545 ;
        RECT 0.000 2485.955 3588.000 2557.745 ;
        RECT 0.000 2481.155 4.160 2485.955 ;
        RECT 3583.840 2481.155 3588.000 2485.955 ;
        RECT 0.000 2409.365 3588.000 2481.155 ;
        RECT 0.000 2404.565 4.160 2409.365 ;
        RECT 3583.840 2404.565 3588.000 2409.365 ;
        RECT 0.000 2332.775 3588.000 2404.565 ;
        RECT 0.000 2327.975 4.160 2332.775 ;
        RECT 3583.840 2327.975 3588.000 2332.775 ;
        RECT 0.000 2256.185 3588.000 2327.975 ;
        RECT 0.000 2251.385 4.160 2256.185 ;
        RECT 3583.840 2251.385 3588.000 2256.185 ;
        RECT 0.000 2179.595 3588.000 2251.385 ;
        RECT 0.000 2174.795 4.160 2179.595 ;
        RECT 3583.840 2174.795 3588.000 2179.595 ;
        RECT 0.000 2103.005 3588.000 2174.795 ;
        RECT 0.000 2098.205 4.160 2103.005 ;
        RECT 3583.840 2098.205 3588.000 2103.005 ;
        RECT 0.000 2026.415 3588.000 2098.205 ;
        RECT 0.000 2021.615 4.160 2026.415 ;
        RECT 3583.840 2021.615 3588.000 2026.415 ;
        RECT 0.000 1949.825 3588.000 2021.615 ;
        RECT 0.000 1945.025 4.160 1949.825 ;
        RECT 3583.840 1945.025 3588.000 1949.825 ;
        RECT 0.000 1873.235 3588.000 1945.025 ;
        RECT 0.000 1868.435 4.160 1873.235 ;
        RECT 3583.840 1868.435 3588.000 1873.235 ;
        RECT 0.000 1796.645 3588.000 1868.435 ;
        RECT 0.000 1791.845 4.160 1796.645 ;
        RECT 3583.840 1791.845 3588.000 1796.645 ;
        RECT 0.000 1720.055 3588.000 1791.845 ;
        RECT 0.000 1715.255 4.160 1720.055 ;
        RECT 3583.840 1715.255 3588.000 1720.055 ;
        RECT 0.000 1643.465 3588.000 1715.255 ;
        RECT 0.000 1638.665 4.160 1643.465 ;
        RECT 3583.840 1638.665 3588.000 1643.465 ;
        RECT 0.000 1566.875 3588.000 1638.665 ;
        RECT 0.000 1562.075 4.160 1566.875 ;
        RECT 3583.840 1562.075 3588.000 1566.875 ;
        RECT 0.000 1490.285 3588.000 1562.075 ;
        RECT 0.000 1485.485 4.160 1490.285 ;
        RECT 3583.840 1485.485 3588.000 1490.285 ;
        RECT 0.000 1413.695 3588.000 1485.485 ;
        RECT 0.000 1408.895 4.160 1413.695 ;
        RECT 3583.840 1408.895 3588.000 1413.695 ;
        RECT 0.000 1337.105 3588.000 1408.895 ;
        RECT 0.000 1332.305 4.160 1337.105 ;
        RECT 3583.840 1332.305 3588.000 1337.105 ;
        RECT 0.000 1260.515 3588.000 1332.305 ;
        RECT 0.000 1255.715 4.160 1260.515 ;
        RECT 3583.840 1255.715 3588.000 1260.515 ;
        RECT 0.000 1183.925 3588.000 1255.715 ;
        RECT 0.000 1179.125 4.160 1183.925 ;
        RECT 3583.840 1179.125 3588.000 1183.925 ;
        RECT 0.000 1107.335 3588.000 1179.125 ;
        RECT 0.000 1102.535 4.160 1107.335 ;
        RECT 3583.840 1102.535 3588.000 1107.335 ;
        RECT 0.000 1030.745 3588.000 1102.535 ;
        RECT 0.000 1025.945 4.160 1030.745 ;
        RECT 3583.840 1025.945 3588.000 1030.745 ;
        RECT 0.000 954.155 3588.000 1025.945 ;
        RECT 0.000 949.355 4.160 954.155 ;
        RECT 3583.840 949.355 3588.000 954.155 ;
        RECT 0.000 877.565 3588.000 949.355 ;
        RECT 0.000 872.765 4.160 877.565 ;
        RECT 3583.840 872.765 3588.000 877.565 ;
        RECT 0.000 800.975 3588.000 872.765 ;
        RECT 0.000 796.175 4.160 800.975 ;
        RECT 3583.840 796.175 3588.000 800.975 ;
        RECT 0.000 724.385 3588.000 796.175 ;
        RECT 0.000 719.585 4.160 724.385 ;
        RECT 3583.840 719.585 3588.000 724.385 ;
        RECT 0.000 647.795 3588.000 719.585 ;
        RECT 0.000 642.995 4.160 647.795 ;
        RECT 3583.840 642.995 3588.000 647.795 ;
        RECT 0.000 571.205 3588.000 642.995 ;
        RECT 0.000 566.405 4.160 571.205 ;
        RECT 3583.840 566.405 3588.000 571.205 ;
        RECT 0.000 494.615 3588.000 566.405 ;
        RECT 0.000 489.815 4.160 494.615 ;
        RECT 3583.840 489.815 3588.000 494.615 ;
        RECT 0.000 418.025 3588.000 489.815 ;
        RECT 0.000 413.225 4.160 418.025 ;
        RECT 3583.840 413.225 3588.000 418.025 ;
        RECT 0.000 341.435 3588.000 413.225 ;
        RECT 0.000 336.635 4.160 341.435 ;
        RECT 3583.840 336.635 3588.000 341.435 ;
        RECT 0.000 264.845 3588.000 336.635 ;
        RECT 0.000 260.045 4.160 264.845 ;
        RECT 3583.840 260.045 3588.000 264.845 ;
        RECT 0.000 188.255 3588.000 260.045 ;
        RECT 0.000 183.455 4.160 188.255 ;
        RECT 3583.840 183.455 3588.000 188.255 ;
        RECT 0.000 111.665 3588.000 183.455 ;
        RECT 0.000 106.865 4.160 111.665 ;
        RECT 3583.840 106.865 3588.000 111.665 ;
        RECT 0.000 35.075 3588.000 106.865 ;
        RECT 0.000 30.275 4.160 35.075 ;
        RECT 3583.840 30.275 3588.000 35.075 ;
        RECT 0.000 0.000 3588.000 30.275 ;
  END
END vsdPLLSoC
END LIBRARY

