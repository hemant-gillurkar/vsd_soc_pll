magic
tech sky130A
magscale 1 2
timestamp 1613927319
<< metal1 >>
rect 39760 920127 39766 920179
rect 39818 920167 39824 920179
rect 282160 920167 282166 920179
rect 39818 920139 282166 920167
rect 39818 920127 39824 920139
rect 282160 920127 282166 920139
rect 282218 920127 282224 920179
rect 282160 917241 282166 917293
rect 282218 917281 282224 917293
rect 303760 917281 303766 917293
rect 282218 917253 303766 917281
rect 282218 917241 282224 917253
rect 303760 917241 303766 917253
rect 303818 917241 303824 917293
rect 303760 912949 303766 913001
rect 303818 912989 303824 913001
rect 303818 912961 308222 912989
rect 303818 912949 303824 912961
rect 308194 912915 308222 912961
rect 313840 912915 313846 912927
rect 308194 912887 313846 912915
rect 313840 912875 313846 912887
rect 313898 912875 313904 912927
rect 313936 904291 313942 904343
rect 313994 904331 314000 904343
rect 318160 904331 318166 904343
rect 313994 904303 318166 904331
rect 313994 904291 314000 904303
rect 318160 904291 318166 904303
rect 318218 904291 318224 904343
rect 318160 796473 318166 796525
rect 318218 796513 318224 796525
rect 323920 796513 323926 796525
rect 318218 796485 323926 796513
rect 318218 796473 318224 796485
rect 323920 796473 323926 796485
rect 323978 796473 323984 796525
rect 323920 757549 323926 757601
rect 323978 757589 323984 757601
rect 326800 757589 326806 757601
rect 323978 757561 326806 757589
rect 323978 757549 323984 757561
rect 326800 757549 326806 757561
rect 326858 757549 326864 757601
rect 326800 665197 326806 665249
rect 326858 665237 326864 665249
rect 329776 665237 329782 665249
rect 326858 665209 329782 665237
rect 326858 665197 326864 665209
rect 329776 665197 329782 665209
rect 329834 665197 329840 665249
rect 329776 651729 329782 651781
rect 329834 651769 329840 651781
rect 332560 651769 332566 651781
rect 329834 651741 332566 651769
rect 329834 651729 329840 651741
rect 332560 651729 332566 651741
rect 332618 651729 332624 651781
rect 332560 615617 332566 615669
rect 332618 615657 332624 615669
rect 334096 615657 334102 615669
rect 332618 615629 334102 615657
rect 332618 615617 332624 615629
rect 334096 615617 334102 615629
rect 334154 615617 334160 615669
rect 334096 601927 334102 601979
rect 334154 601967 334160 601979
rect 339856 601967 339862 601979
rect 334154 601939 339862 601967
rect 334154 601927 334160 601939
rect 339856 601927 339862 601939
rect 339914 601927 339920 601979
rect 345904 518603 345910 518655
rect 345962 518643 345968 518655
rect 625840 518643 625846 518655
rect 345962 518615 625846 518643
rect 345962 518603 345968 518615
rect 625840 518603 625846 518615
rect 625898 518603 625904 518655
rect 329680 511203 329686 511255
rect 329738 511243 329744 511255
rect 347056 511243 347062 511255
rect 329738 511215 347062 511243
rect 329738 511203 329744 511215
rect 347056 511203 347062 511215
rect 347114 511203 347120 511255
rect 625840 508761 625846 508813
rect 625898 508801 625904 508813
rect 629200 508801 629206 508813
rect 625898 508773 629206 508801
rect 625898 508761 625904 508773
rect 629200 508761 629206 508773
rect 629258 508761 629264 508813
rect 317968 495367 317974 495419
rect 318026 495407 318032 495419
rect 329680 495407 329686 495419
rect 318026 495379 329686 495407
rect 318026 495367 318032 495379
rect 329680 495367 329686 495379
rect 329738 495367 329744 495419
rect 306640 485155 306646 485207
rect 306698 485195 306704 485207
rect 317968 485195 317974 485207
rect 306698 485167 317974 485195
rect 306698 485155 306704 485167
rect 317968 485155 317974 485167
rect 318026 485155 318032 485207
rect 629200 474573 629206 474625
rect 629258 474613 629264 474625
rect 632176 474613 632182 474625
rect 629258 474585 632182 474613
rect 629258 474573 629264 474585
rect 632176 474573 632182 474585
rect 632234 474573 632240 474625
rect 39856 472279 39862 472331
rect 39914 472319 39920 472331
rect 306640 472319 306646 472331
rect 39914 472291 306646 472319
rect 39914 472279 39920 472291
rect 306640 472279 306646 472291
rect 306698 472279 306704 472331
rect 632176 469393 632182 469445
rect 632234 469433 632240 469445
rect 634960 469433 634966 469445
rect 632234 469405 634966 469433
rect 632234 469393 632240 469405
rect 634960 469393 634966 469405
rect 635018 469393 635024 469445
rect 634960 411747 634966 411799
rect 635018 411787 635024 411799
rect 636496 411787 636502 411799
rect 635018 411759 636502 411787
rect 635018 411747 635024 411759
rect 636496 411747 636502 411759
rect 636554 411747 636560 411799
rect 636496 408861 636502 408913
rect 636554 408901 636560 408913
rect 640240 408901 640246 408913
rect 636554 408873 640246 408901
rect 636554 408861 636560 408873
rect 640240 408861 640246 408873
rect 640298 408861 640304 408913
rect 640240 400277 640246 400329
rect 640298 400317 640304 400329
rect 643600 400317 643606 400329
rect 640298 400289 643606 400317
rect 640298 400277 640304 400289
rect 643600 400277 643606 400289
rect 643658 400277 643664 400329
rect 498256 391693 498262 391745
rect 498314 391733 498320 391745
rect 675018 391733 675024 391745
rect 498314 391705 675024 391733
rect 498314 391693 498320 391705
rect 675018 391693 675024 391705
rect 675076 391693 675082 391745
rect 643600 359947 643606 359999
rect 643658 359987 643664 359999
rect 653776 359987 653782 359999
rect 643658 359959 653782 359987
rect 643658 359947 643664 359959
rect 653776 359947 653782 359959
rect 653834 359947 653840 359999
rect 653776 357061 653782 357113
rect 653834 357101 653840 357113
rect 660880 357101 660886 357113
rect 653834 357073 660886 357101
rect 653834 357061 653840 357073
rect 660880 357061 660886 357073
rect 660938 357061 660944 357113
rect 660880 319617 660886 319669
rect 660938 319657 660944 319669
rect 663760 319657 663766 319669
rect 660938 319629 663766 319657
rect 660938 319617 660944 319629
rect 663760 319617 663766 319629
rect 663818 319617 663824 319669
rect 498256 307925 498262 307977
rect 498314 307965 498320 307977
rect 500368 307965 500374 307977
rect 498314 307937 500374 307965
rect 498314 307925 498320 307937
rect 500368 307925 500374 307937
rect 500426 307925 500432 307977
rect 663760 293865 663766 293917
rect 663818 293905 663824 293917
rect 666640 293905 666646 293917
rect 663818 293877 666646 293905
rect 663818 293865 663824 293877
rect 666640 293865 666646 293877
rect 666698 293865 666704 293917
rect 666640 275513 666646 275565
rect 666698 275553 666704 275565
rect 669616 275553 669622 275565
rect 666698 275525 669622 275553
rect 666698 275513 666704 275525
rect 669616 275513 669622 275525
rect 669674 275513 669680 275565
rect 669616 262045 669622 262097
rect 669674 262085 669680 262097
rect 672400 262085 672406 262097
rect 669674 262057 672406 262085
rect 669674 262045 669680 262057
rect 672400 262045 672406 262057
rect 672458 262045 672464 262097
rect 672400 241843 672406 241895
rect 672458 241883 672464 241895
rect 675280 241883 675286 241895
rect 672458 241855 675286 241883
rect 672458 241843 672464 241855
rect 675280 241843 675286 241855
rect 675338 241843 675344 241895
rect 675280 215129 675286 215181
rect 675338 215169 675344 215181
rect 677104 215169 677110 215181
rect 675338 215141 677110 215169
rect 675338 215129 675344 215141
rect 677104 215129 677110 215141
rect 677162 215129 677168 215181
rect 677104 213057 677110 213109
rect 677162 213097 677168 213109
rect 682480 213097 682486 213109
rect 677162 213069 682486 213097
rect 677162 213057 677168 213069
rect 682480 213057 682486 213069
rect 682538 213057 682544 213109
rect 682576 201587 682582 201639
rect 682634 201627 682640 201639
rect 682634 201599 694142 201627
rect 682634 201587 682640 201599
rect 694114 201553 694142 201599
rect 699760 201553 699766 201565
rect 694114 201525 699766 201553
rect 699760 201513 699766 201525
rect 699818 201513 699824 201565
<< via1 >>
rect 39766 920127 39818 920179
rect 282166 920127 282218 920179
rect 282166 917241 282218 917293
rect 303766 917241 303818 917293
rect 303766 912949 303818 913001
rect 313846 912875 313898 912927
rect 313942 904291 313994 904343
rect 318166 904291 318218 904343
rect 318166 796473 318218 796525
rect 323926 796473 323978 796525
rect 323926 757549 323978 757601
rect 326806 757549 326858 757601
rect 326806 665197 326858 665249
rect 329782 665197 329834 665249
rect 329782 651729 329834 651781
rect 332566 651729 332618 651781
rect 332566 615617 332618 615669
rect 334102 615617 334154 615669
rect 334102 601927 334154 601979
rect 339862 601927 339914 601979
rect 345910 518603 345962 518655
rect 625846 518603 625898 518655
rect 329686 511203 329738 511255
rect 347062 511203 347114 511255
rect 625846 508761 625898 508813
rect 629206 508761 629258 508813
rect 317974 495367 318026 495419
rect 329686 495367 329738 495419
rect 306646 485155 306698 485207
rect 317974 485155 318026 485207
rect 629206 474573 629258 474625
rect 632182 474573 632234 474625
rect 39862 472279 39914 472331
rect 306646 472279 306698 472331
rect 632182 469393 632234 469445
rect 634966 469393 635018 469445
rect 634966 411747 635018 411799
rect 636502 411747 636554 411799
rect 636502 408861 636554 408913
rect 640246 408861 640298 408913
rect 640246 400277 640298 400329
rect 643606 400277 643658 400329
rect 498262 391693 498314 391745
rect 675024 391693 675076 391745
rect 643606 359947 643658 359999
rect 653782 359947 653834 359999
rect 653782 357061 653834 357113
rect 660886 357061 660938 357113
rect 660886 319617 660938 319669
rect 663766 319617 663818 319669
rect 498262 307925 498314 307977
rect 500374 307925 500426 307977
rect 663766 293865 663818 293917
rect 666646 293865 666698 293917
rect 666646 275513 666698 275565
rect 669622 275513 669674 275565
rect 669622 262045 669674 262097
rect 672406 262045 672458 262097
rect 672406 241843 672458 241895
rect 675286 241843 675338 241895
rect 675286 215129 675338 215181
rect 677110 215129 677162 215181
rect 677110 213057 677162 213109
rect 682486 213057 682538 213109
rect 682582 201587 682634 201639
rect 699766 201513 699818 201565
<< metal2 >>
rect 39764 920218 39820 920227
rect 39764 920153 39766 920162
rect 39818 920153 39820 920162
rect 282166 920179 282218 920185
rect 39766 920121 39818 920127
rect 282166 920121 282218 920127
rect 282178 917299 282206 920121
rect 282166 917293 282218 917299
rect 282166 917235 282218 917241
rect 303766 917293 303818 917299
rect 303766 917235 303818 917241
rect 303778 913007 303806 917235
rect 303766 913001 303818 913007
rect 303766 912943 303818 912949
rect 313846 912927 313898 912933
rect 313846 912869 313898 912875
rect 313858 907180 313886 912869
rect 313858 907152 313982 907180
rect 313954 904349 313982 907152
rect 313942 904343 313994 904349
rect 313942 904285 313994 904291
rect 318166 904343 318218 904349
rect 318166 904285 318218 904291
rect 42178 835275 42206 835645
rect 42164 835266 42220 835275
rect 42164 835201 42220 835210
rect 318178 796531 318206 904285
rect 318166 796525 318218 796531
rect 318166 796467 318218 796473
rect 323926 796525 323978 796531
rect 323926 796467 323978 796473
rect 323938 757607 323966 796467
rect 323926 757601 323978 757607
rect 323926 757543 323978 757549
rect 326806 757601 326858 757607
rect 326806 757543 326858 757549
rect 42178 746179 42206 746660
rect 42164 746170 42220 746179
rect 42164 746105 42220 746114
rect 326818 665255 326846 757543
rect 326806 665249 326858 665255
rect 326806 665191 326858 665197
rect 329782 665249 329834 665255
rect 329782 665191 329834 665197
rect 329794 651787 329822 665191
rect 329782 651781 329834 651787
rect 329782 651723 329834 651729
rect 332566 651781 332618 651787
rect 332566 651723 332618 651729
rect 332578 615675 332606 651723
rect 332566 615669 332618 615675
rect 332566 615611 332618 615617
rect 334102 615669 334154 615675
rect 334102 615611 334154 615617
rect 334114 601985 334142 615611
rect 334102 601979 334154 601985
rect 334102 601921 334154 601927
rect 339862 601979 339914 601985
rect 339862 601921 339914 601927
rect 339874 520479 339902 601921
rect 340628 520914 340684 520923
rect 340628 520849 340684 520858
rect 339860 520470 339916 520479
rect 339860 520405 339916 520414
rect 340642 519998 340670 520849
rect 340820 519878 340876 519887
rect 340820 519813 340876 519822
rect 340834 519406 340862 519813
rect 345910 518655 345962 518661
rect 345910 518597 345962 518603
rect 345922 518370 345950 518597
rect 347074 511261 347102 519702
rect 625846 518655 625898 518661
rect 625846 518597 625898 518603
rect 329686 511255 329738 511261
rect 329686 511197 329738 511203
rect 347062 511255 347114 511261
rect 347062 511197 347114 511203
rect 329698 495425 329726 511197
rect 625858 508819 625886 518597
rect 625846 508813 625898 508819
rect 625846 508755 625898 508761
rect 629206 508813 629258 508819
rect 629206 508755 629258 508761
rect 317974 495419 318026 495425
rect 317974 495361 318026 495367
rect 329686 495419 329738 495425
rect 329686 495361 329738 495367
rect 317986 485213 318014 495361
rect 306646 485207 306698 485213
rect 306646 485149 306698 485155
rect 317974 485207 318026 485213
rect 317974 485149 318026 485155
rect 39860 476070 39916 476079
rect 39860 476005 39916 476014
rect 39874 472337 39902 476005
rect 306658 472337 306686 485149
rect 629218 474631 629246 508755
rect 629206 474625 629258 474631
rect 629206 474567 629258 474573
rect 632182 474625 632234 474631
rect 632182 474567 632234 474573
rect 39862 472331 39914 472337
rect 39862 472273 39914 472279
rect 306646 472331 306698 472337
rect 306646 472273 306698 472279
rect 632194 469451 632222 474567
rect 632182 469445 632234 469451
rect 632182 469387 632234 469393
rect 634966 469445 635018 469451
rect 634966 469387 635018 469393
rect 634978 411805 635006 469387
rect 634966 411799 635018 411805
rect 634966 411741 635018 411747
rect 636502 411799 636554 411805
rect 636502 411741 636554 411747
rect 636514 408919 636542 411741
rect 636502 408913 636554 408919
rect 636502 408855 636554 408861
rect 640246 408913 640298 408919
rect 640246 408855 640298 408861
rect 640258 400335 640286 408855
rect 640246 400329 640298 400335
rect 640246 400271 640298 400277
rect 643606 400329 643658 400335
rect 643606 400271 643658 400277
rect 498262 391745 498314 391751
rect 498262 391687 498314 391693
rect 498274 307983 498302 391687
rect 643618 360005 643646 400271
rect 675024 391745 675076 391751
rect 675024 391687 675076 391693
rect 675036 391682 675064 391687
rect 643606 359999 643658 360005
rect 643606 359941 643658 359947
rect 653782 359999 653834 360005
rect 653782 359941 653834 359947
rect 653794 357119 653822 359941
rect 653782 357113 653834 357119
rect 653782 357055 653834 357061
rect 660886 357113 660938 357119
rect 660886 357055 660938 357061
rect 660898 319675 660926 357055
rect 660886 319669 660938 319675
rect 660886 319611 660938 319617
rect 663766 319669 663818 319675
rect 663766 319611 663818 319617
rect 498262 307977 498314 307983
rect 498262 307919 498314 307925
rect 500374 307977 500426 307983
rect 500374 307919 500426 307925
rect 500386 299788 500414 307919
rect 500386 299760 500784 299788
rect 663778 293923 663806 319611
rect 663766 293917 663818 293923
rect 663766 293859 663818 293865
rect 666646 293917 666698 293923
rect 666646 293859 666698 293865
rect 666658 275571 666686 293859
rect 666646 275565 666698 275571
rect 666646 275507 666698 275513
rect 669622 275565 669674 275571
rect 669622 275507 669674 275513
rect 669634 262103 669662 275507
rect 669622 262097 669674 262103
rect 669622 262039 669674 262045
rect 672406 262097 672458 262103
rect 672406 262039 672458 262045
rect 672418 241901 672446 262039
rect 672406 241895 672458 241901
rect 672406 241837 672458 241843
rect 675286 241895 675338 241901
rect 675286 241837 675338 241843
rect 675298 215187 675326 241837
rect 675286 215181 675338 215187
rect 675286 215123 675338 215129
rect 677110 215181 677162 215187
rect 677110 215123 677162 215129
rect 677122 213115 677150 215123
rect 677110 213109 677162 213115
rect 677110 213051 677162 213057
rect 682486 213109 682538 213115
rect 682486 213051 682538 213057
rect 682498 207288 682526 213051
rect 682498 207260 682622 207288
rect 682594 201645 682622 207260
rect 682582 201639 682634 201645
rect 682582 201581 682634 201587
rect 699766 201565 699818 201571
rect 699766 201507 699818 201513
rect 699778 192932 699806 201507
rect 699778 192904 699902 192932
rect 699874 161135 699902 192904
rect 677780 161126 677836 161135
rect 677780 161061 677836 161070
rect 699860 161126 699916 161135
rect 699860 161061 699916 161070
rect 677794 150651 677822 161061
rect 677780 150642 677836 150651
rect 677780 150577 677836 150586
<< via2 >>
rect 39764 920179 39820 920218
rect 39764 920162 39766 920179
rect 39766 920162 39818 920179
rect 39818 920162 39820 920179
rect 42164 835210 42220 835266
rect 42164 746114 42220 746170
rect 340628 520858 340684 520914
rect 339860 520414 339916 520470
rect 340820 519822 340876 519878
rect 39860 476014 39916 476070
rect 677780 161070 677836 161126
rect 699860 161070 699916 161126
rect 677780 150586 677836 150642
<< metal3 >>
rect 39759 920220 39825 920223
rect 39456 920218 39825 920220
rect 39456 920162 39764 920218
rect 39820 920162 39825 920218
rect 39456 920160 39825 920162
rect 39759 920157 39825 920160
rect 42159 835268 42225 835271
rect 43066 835268 43072 835270
rect 42159 835266 43072 835268
rect 42159 835210 42164 835266
rect 42220 835210 43072 835266
rect 42159 835208 43072 835210
rect 42159 835205 42225 835208
rect 43066 835206 43072 835208
rect 43136 835206 43142 835270
rect 42159 746172 42225 746175
rect 42874 746172 42880 746174
rect 42159 746170 42880 746172
rect 42159 746114 42164 746170
rect 42220 746114 42880 746170
rect 42159 746112 42880 746114
rect 42159 746109 42225 746112
rect 42874 746110 42880 746112
rect 42944 746110 42950 746174
rect 42874 520854 42880 520918
rect 42944 520916 42950 520918
rect 340623 520916 340689 520919
rect 42944 520914 340689 520916
rect 42944 520858 340628 520914
rect 340684 520858 340689 520914
rect 42944 520856 340689 520858
rect 42944 520854 42950 520856
rect 340623 520853 340689 520856
rect 43066 520706 43072 520770
rect 43136 520768 43142 520770
rect 43136 520708 338814 520768
rect 43136 520706 43142 520708
rect 338754 520324 338814 520708
rect 339855 520472 339921 520475
rect 339855 520470 341472 520472
rect 339855 520414 339860 520470
rect 339916 520414 341472 520470
rect 339855 520412 341472 520414
rect 339855 520409 339921 520412
rect 338754 520264 340926 520324
rect 340866 519883 340926 520264
rect 340815 519878 340926 519883
rect 340815 519822 340820 519878
rect 340876 519822 340926 519878
rect 340815 519820 340926 519822
rect 340815 519817 340881 519820
rect 39855 476072 39921 476075
rect 25824 476070 39921 476072
rect 25824 476014 39860 476070
rect 39916 476014 39921 476070
rect 25824 476012 39921 476014
rect 39855 476009 39921 476012
rect 677775 161128 677841 161131
rect 699855 161128 699921 161131
rect 677775 161126 699921 161128
rect 677775 161070 677780 161126
rect 677836 161070 699860 161126
rect 699916 161070 699921 161126
rect 677775 161068 699921 161070
rect 677775 161065 677841 161068
rect 699855 161065 699921 161068
rect 677775 150644 677841 150647
rect 677775 150642 678048 150644
rect 677775 150586 677780 150642
rect 677836 150586 678048 150642
rect 677775 150584 678048 150586
rect 677775 150581 677841 150584
<< via3 >>
rect 43072 835206 43136 835270
rect 42880 746110 42944 746174
rect 42880 520854 42944 520918
rect 43072 520706 43136 520770
<< metal4 >>
rect 43071 835270 43137 835271
rect 43071 835206 43072 835270
rect 43136 835206 43137 835270
rect 43071 835205 43137 835206
rect 42879 746174 42945 746175
rect 42879 746110 42880 746174
rect 42944 746110 42945 746174
rect 42879 746109 42945 746110
rect 42882 520919 42942 746109
rect 42879 520918 42945 520919
rect 42879 520854 42880 520918
rect 42944 520854 42945 520918
rect 42879 520853 42945 520854
rect 43074 520771 43134 835205
rect 43071 520770 43137 520771
rect 43071 520706 43072 520770
rect 43136 520706 43137 520770
rect 43071 520705 43137 520706
<< metal5 >>
rect 1152 1032681 716448 1033001
rect 1152 1017363 716448 1017683
rect 1152 1002045 716448 1002365
rect 1152 986727 716448 987047
rect 1152 971409 716448 971729
rect 1152 956091 716448 956411
rect 1152 940773 716448 941093
rect 1152 925455 716448 925775
rect 1152 910137 716448 910457
rect 1152 894819 716448 895139
rect 1152 879501 716448 879821
rect 1152 864183 716448 864503
rect 1152 848865 716448 849185
rect 1152 833547 716448 833867
rect 1152 818229 716448 818549
rect 1152 802911 716448 803231
rect 1152 787593 716448 787913
rect 1152 772275 716448 772595
rect 1152 756957 716448 757277
rect 1152 741639 716448 741959
rect 1152 726321 716448 726641
rect 1152 711003 716448 711323
rect 1152 695685 716448 696005
rect 1152 680367 716448 680687
rect 1152 665049 716448 665369
rect 1152 649731 716448 650051
rect 1152 634413 716448 634733
rect 1152 619095 716448 619415
rect 1152 603777 716448 604097
rect 1152 588459 716448 588779
rect 1152 573141 716448 573461
rect 1152 557823 716448 558143
rect 1152 542505 716448 542825
rect 1152 527187 716448 527507
rect 1152 511869 716448 512189
rect 1152 496551 716448 496871
rect 1152 481233 716448 481553
rect 1152 465915 716448 466235
rect 1152 450597 716448 450917
rect 1152 435279 716448 435599
rect 1152 419961 716448 420281
rect 1152 404643 716448 404963
rect 1152 389325 716448 389645
rect 1152 374007 716448 374327
rect 1152 358689 716448 359009
rect 1152 343371 716448 343691
rect 1152 328053 716448 328373
rect 1152 312735 716448 313055
rect 1152 297417 716448 297737
rect 1152 282099 716448 282419
rect 1152 266781 716448 267101
rect 1152 251463 716448 251783
rect 1152 236145 716448 236465
rect 1152 220827 716448 221147
rect 1152 205509 716448 205829
rect 1152 190191 716448 190511
rect 1152 174873 716448 175193
rect 1152 159555 716448 159875
rect 1152 144237 716448 144557
rect 1152 128919 716448 129239
rect 1152 113601 716448 113921
rect 1152 98283 716448 98603
rect 1152 82965 716448 83285
rect 1152 67647 716448 67967
rect 1152 52329 716448 52649
rect 1152 37011 716448 37331
rect 1152 21693 716448 22013
rect 1152 6375 716448 6695
use simple_por  POR
timestamp 1613927319
transform 1 0 500000 0 -1 308164
box 0 0 4360 9164
use avsdpll_1v8  PLL
timestamp 1613927319
transform 1 0 340000 0 1 518000
box 0 0 7236 2742
use chip_io  PADFRAME
timestamp 1613927319
transform 1 0 0 0 1 0
box 0 0 717600 1037600
<< labels >>
rlabel metal5 s 1152 1017363 716448 1017683 6 VPWR
port 0 nsew power bidirectional
rlabel metal5 s 1152 986727 716448 987047 6 VPWR.extra1
port 1 nsew power bidirectional
rlabel metal5 s 1152 956091 716448 956411 6 VPWR.extra2
port 2 nsew power bidirectional
rlabel metal5 s 1152 925455 716448 925775 6 VPWR.extra3
port 3 nsew power bidirectional
rlabel metal5 s 1152 894819 716448 895139 6 VPWR.extra4
port 4 nsew power bidirectional
rlabel metal5 s 1152 864183 716448 864503 6 VPWR.extra5
port 5 nsew power bidirectional
rlabel metal5 s 1152 833547 716448 833867 6 VPWR.extra6
port 6 nsew power bidirectional
rlabel metal5 s 1152 802911 716448 803231 6 VPWR.extra7
port 7 nsew power bidirectional
rlabel metal5 s 1152 772275 716448 772595 6 VPWR.extra8
port 8 nsew power bidirectional
rlabel metal5 s 1152 741639 716448 741959 6 VPWR.extra9
port 9 nsew power bidirectional
rlabel metal5 s 1152 711003 716448 711323 6 VPWR.extra10
port 10 nsew power bidirectional
rlabel metal5 s 1152 680367 716448 680687 6 VPWR.extra11
port 11 nsew power bidirectional
rlabel metal5 s 1152 649731 716448 650051 6 VPWR.extra12
port 12 nsew power bidirectional
rlabel metal5 s 1152 619095 716448 619415 6 VPWR.extra13
port 13 nsew power bidirectional
rlabel metal5 s 1152 588459 716448 588779 6 VPWR.extra14
port 14 nsew power bidirectional
rlabel metal5 s 1152 557823 716448 558143 6 VPWR.extra15
port 15 nsew power bidirectional
rlabel metal5 s 1152 527187 716448 527507 6 VPWR.extra16
port 16 nsew power bidirectional
rlabel metal5 s 1152 496551 716448 496871 6 VPWR.extra17
port 17 nsew power bidirectional
rlabel metal5 s 1152 465915 716448 466235 6 VPWR.extra18
port 18 nsew power bidirectional
rlabel metal5 s 1152 435279 716448 435599 6 VPWR.extra19
port 19 nsew power bidirectional
rlabel metal5 s 1152 404643 716448 404963 6 VPWR.extra20
port 20 nsew power bidirectional
rlabel metal5 s 1152 374007 716448 374327 6 VPWR.extra21
port 21 nsew power bidirectional
rlabel metal5 s 1152 343371 716448 343691 6 VPWR.extra22
port 22 nsew power bidirectional
rlabel metal5 s 1152 312735 716448 313055 6 VPWR.extra23
port 23 nsew power bidirectional
rlabel metal5 s 1152 282099 716448 282419 6 VPWR.extra24
port 24 nsew power bidirectional
rlabel metal5 s 1152 251463 716448 251783 6 VPWR.extra25
port 25 nsew power bidirectional
rlabel metal5 s 1152 220827 716448 221147 6 VPWR.extra26
port 26 nsew power bidirectional
rlabel metal5 s 1152 190191 716448 190511 6 VPWR.extra27
port 27 nsew power bidirectional
rlabel metal5 s 1152 159555 716448 159875 6 VPWR.extra28
port 28 nsew power bidirectional
rlabel metal5 s 1152 128919 716448 129239 6 VPWR.extra29
port 29 nsew power bidirectional
rlabel metal5 s 1152 98283 716448 98603 6 VPWR.extra30
port 30 nsew power bidirectional
rlabel metal5 s 1152 67647 716448 67967 6 VPWR.extra31
port 31 nsew power bidirectional
rlabel metal5 s 1152 37011 716448 37331 6 VPWR.extra32
port 32 nsew power bidirectional
rlabel metal5 s 1152 6375 716448 6695 6 VPWR.extra33
port 33 nsew power bidirectional
rlabel metal5 s 1152 1032681 716448 1033001 6 VGND
port 34 nsew ground bidirectional
rlabel metal5 s 1152 1002045 716448 1002365 6 VGND.extra1
port 35 nsew ground bidirectional
rlabel metal5 s 1152 971409 716448 971729 6 VGND.extra2
port 36 nsew ground bidirectional
rlabel metal5 s 1152 940773 716448 941093 6 VGND.extra3
port 37 nsew ground bidirectional
rlabel metal5 s 1152 910137 716448 910457 6 VGND.extra4
port 38 nsew ground bidirectional
rlabel metal5 s 1152 879501 716448 879821 6 VGND.extra5
port 39 nsew ground bidirectional
rlabel metal5 s 1152 848865 716448 849185 6 VGND.extra6
port 40 nsew ground bidirectional
rlabel metal5 s 1152 818229 716448 818549 6 VGND.extra7
port 41 nsew ground bidirectional
rlabel metal5 s 1152 787593 716448 787913 6 VGND.extra8
port 42 nsew ground bidirectional
rlabel metal5 s 1152 756957 716448 757277 6 VGND.extra9
port 43 nsew ground bidirectional
rlabel metal5 s 1152 726321 716448 726641 6 VGND.extra10
port 44 nsew ground bidirectional
rlabel metal5 s 1152 695685 716448 696005 6 VGND.extra11
port 45 nsew ground bidirectional
rlabel metal5 s 1152 665049 716448 665369 6 VGND.extra12
port 46 nsew ground bidirectional
rlabel metal5 s 1152 634413 716448 634733 6 VGND.extra13
port 47 nsew ground bidirectional
rlabel metal5 s 1152 603777 716448 604097 6 VGND.extra14
port 48 nsew ground bidirectional
rlabel metal5 s 1152 573141 716448 573461 6 VGND.extra15
port 49 nsew ground bidirectional
rlabel metal5 s 1152 542505 716448 542825 6 VGND.extra16
port 50 nsew ground bidirectional
rlabel metal5 s 1152 511869 716448 512189 6 VGND.extra17
port 51 nsew ground bidirectional
rlabel metal5 s 1152 481233 716448 481553 6 VGND.extra18
port 52 nsew ground bidirectional
rlabel metal5 s 1152 450597 716448 450917 6 VGND.extra19
port 53 nsew ground bidirectional
rlabel metal5 s 1152 419961 716448 420281 6 VGND.extra20
port 54 nsew ground bidirectional
rlabel metal5 s 1152 389325 716448 389645 6 VGND.extra21
port 55 nsew ground bidirectional
rlabel metal5 s 1152 358689 716448 359009 6 VGND.extra22
port 56 nsew ground bidirectional
rlabel metal5 s 1152 328053 716448 328373 6 VGND.extra23
port 57 nsew ground bidirectional
rlabel metal5 s 1152 297417 716448 297737 6 VGND.extra24
port 58 nsew ground bidirectional
rlabel metal5 s 1152 266781 716448 267101 6 VGND.extra25
port 59 nsew ground bidirectional
rlabel metal5 s 1152 236145 716448 236465 6 VGND.extra26
port 60 nsew ground bidirectional
rlabel metal5 s 1152 205509 716448 205829 6 VGND.extra27
port 61 nsew ground bidirectional
rlabel metal5 s 1152 174873 716448 175193 6 VGND.extra28
port 62 nsew ground bidirectional
rlabel metal5 s 1152 144237 716448 144557 6 VGND.extra29
port 63 nsew ground bidirectional
rlabel metal5 s 1152 113601 716448 113921 6 VGND.extra30
port 64 nsew ground bidirectional
rlabel metal5 s 1152 82965 716448 83285 6 VGND.extra31
port 65 nsew ground bidirectional
rlabel metal5 s 1152 52329 716448 52649 6 VGND.extra32
port 66 nsew ground bidirectional
rlabel metal5 s 1152 21693 716448 22013 6 VGND.extra33
port 67 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 717600 1037600
<< end >>
